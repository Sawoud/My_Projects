/*
Copyright by Henry Ko and Nicola Nicolici
Department of Electrical and Computer Engineering
McMaster University
Ontario, Canada
*/

`timescale 1ns/100ps
`ifndef DISABLE_DEFAULT_NET
`default_nettype none
`endif

`include "define_state.h"

// This is the top module
// It connects the UART, SRAM and VGA together.
// It gives access to the SRAM for UART and VGA
module experiment4 (
		/////// board clocks                      ////////////
		input logic CLOCK_50_I,                   // 50 MHz clock

		/////// pushbuttons/switches              ////////////
		input logic[3:0] PUSH_BUTTON_N_I,         // pushbuttons
		input logic[17:0] SWITCH_I,               // toggle switches

		/////// 7 segment displays/LEDs           ////////////
		output logic[6:0] SEVEN_SEGMENT_N_O[7:0], // 8 seven segment displays
		output logic[8:0] LED_GREEN_O,            // 9 green LEDs

		/////// VGA interface                     ////////////
		output logic VGA_CLOCK_O,                 // VGA clock
		output logic VGA_HSYNC_O,                 // VGA H_SYNC
		output logic VGA_VSYNC_O,                 // VGA V_SYNC
		output logic VGA_BLANK_O,                 // VGA BLANK
		output logic VGA_SYNC_O,                  // VGA SYNC
		output logic[7:0] VGA_RED_O,              // VGA red
		output logic[7:0] VGA_GREEN_O,            // VGA green
		output logic[7:0] VGA_BLUE_O,             // VGA blue
		
		/////// SRAM Interface                    ////////////
		inout wire[15:0] SRAM_DATA_IO,            // SRAM data bus 16 bits
		output logic[19:0] SRAM_ADDRESS_O,        // SRAM address bus 18 bits
		output logic SRAM_UB_N_O,                 // SRAM high-byte data mask 
		output logic SRAM_LB_N_O,                 // SRAM low-byte data mask 
		output logic SRAM_WE_N_O,                 // SRAM write enable
		output logic SRAM_CE_N_O,                 // SRAM chip enable
		output logic SRAM_OE_N_O,                 // SRAM output logic enable
		
		/////// UART                              ////////////
		input  logic UART_RX_I,                   // UART receive signal
		output logic UART_TX_O                    // UART transmit signal
);
	
logic resetn;

upsample_type upsample;

// For M1
logic [17:0] M1_Address;
logic [15:0] M1_write_data;
logic [31:0] Up [76799:0];
logic [31:0] Up [76799:0];

logic M1_wr_n, M1_start, M1_finish;

// For Push button
logic [3:0] PB_pushed;

// For VGA SRAM interface
logic VGA_enable;
logic [17:0] VGA_base_address;
logic [17:0] VGA_SRAM_address;

// For SRAM
logic [17:0] SRAM_address;
logic [15:0] SRAM_write_data;
logic SRAM_we_n;
logic [15:0] SRAM_read_data;
logic SRAM_ready;

// For UART SRAM interface
logic UART_rx_enable;
logic UART_rx_initialize;
logic [17:0] UART_SRAM_address;
logic [15:0] UART_SRAM_write_data;
logic UART_SRAM_we_n;
logic [25:0] UART_timer;

logic [6:0] value_7_segment [7:0];

// For error detection in UART
logic Frame_error;

// For disabling UART transmit
assign UART_TX_O = 1'b1;

assign resetn = ~SWITCH_I[17] && SRAM_ready;

// M1 Module
M1 M1_interface (
	.Clock(CLOCK_50_I),
	.Resetn(resetn),
	.SRAM_read_data(SRAM_read_data),
	.M1_Address(M1_Address),
	.M1_write_data(M1_write_data),
	.M1_wr_n(M1_wr_n),
	.M1_start(M1_start),
	.M1_finish(M1_finish)
);

// Push Button unit
PB_controller PB_unit (
	.Clock_50(CLOCK_50_I),
	.Resetn(resetn),
	.PB_signal(PUSH_BUTTON_N_I),	
	.PB_pushed(PB_pushed)
);

VGA_SRAM_interface VGA_unit (
	.Clock(CLOCK_50_I),
	.Resetn(resetn),
	.VGA_enable(VGA_enable),
   
	// For accessing SRAM
	.SRAM_base_address(VGA_base_address),
	.SRAM_address(VGA_SRAM_address),
	.SRAM_read_data(SRAM_read_data),
   
	// To VGA pins
	.VGA_CLOCK_O(VGA_CLOCK_O),
	.VGA_HSYNC_O(VGA_HSYNC_O),
	.VGA_VSYNC_O(VGA_VSYNC_O),
	.VGA_BLANK_O(VGA_BLANK_O),
	.VGA_SYNC_O(VGA_SYNC_O),
	.VGA_RED_O(VGA_RED_O),
	.VGA_GREEN_O(VGA_GREEN_O),
	.VGA_BLUE_O(VGA_BLUE_O)
);

// UART SRAM interface
UART_SRAM_interface UART_unit(
	.Clock(CLOCK_50_I),
	.Resetn(resetn), 
   
	.UART_RX_I(UART_RX_I),
	.Initialize(UART_rx_initialize),
	.Enable(UART_rx_enable),
   
	// For accessing SRAM
	.SRAM_address(UART_SRAM_address),
	.SRAM_write_data(UART_SRAM_write_data),
	.SRAM_we_n(UART_SRAM_we_n),
	.Frame_error(Frame_error)
);

// SRAM unit
SRAM_controller SRAM_unit (
	.Clock_50(CLOCK_50_I),
	.Resetn(~SWITCH_I[17]),
	.SRAM_address(SRAM_address),
	.SRAM_write_data(SRAM_write_data),
	.SRAM_we_n(SRAM_we_n),
	.SRAM_read_data(SRAM_read_data),		
	.SRAM_ready(SRAM_ready),
		
	// To the SRAM pins
	.SRAM_DATA_IO(SRAM_DATA_IO),
	.SRAM_ADDRESS_O(SRAM_ADDRESS_O[17:0]),
	.SRAM_UB_N_O(SRAM_UB_N_O),
	.SRAM_LB_N_O(SRAM_LB_N_O),
	.SRAM_WE_N_O(SRAM_WE_N_O),
	.SRAM_CE_N_O(SRAM_CE_N_O),
	.SRAM_OE_N_O(SRAM_OE_N_O)
);
logic [15:0] Ru [5:0];
logic [15:0] Rv [5:0];
logic [31:0] ACC [4:0];

logic MULT1_IN_1[31:0];
logic MULT1_IN_2[31:0];
logic MULT1_OUT_1 [63:0];

logic MULT2_IN_1[31:0];
logic MULT2_IN_2[31:0];
logic MULT2_OUT_1 [63:0];

logic MULT3_IN_1[31:0];
logic MULT3_IN_2[31:0];
logic MULT3_OUT_1 [63:0];

logic MULT4_IN_1[31:0];
logic MULT4_IN_2[31:0];
logic MULT4_OUT_1 [63:0];

assign SRAM_ADDRESS_O[19:18] = 2'b00;

// Give access to SRAM for UART and VGA at appropriate time
	assign SRAM_address = 16'd38400;

	assign SRAM_write_data = 16'd0;

	assign SRAM_we_n =  1'b1;
	integer j;

always @(posedge CLOCK_50_I or negedge resetn) begin
	if (~resetn) begin
		top_state <= S_IDLE;
		
		UART_rx_initialize <= 1'b0;
		UART_rx_enable <= 1'b0;
		UART_timer <= 26'd0;
		j <= 0;
		VGA_enable <= 1'b1;
		shift_reg[5:0];
		integer i;
	end else begin

		// By default the UART timer (used for timeout detection) is incremented
		// it will be synchronously reset to 0 under a few conditions (see below)

		case (upsample)
		SL0: begin
				Ru[0] = SRAM_read_data[15:8];
				MULT1_IN_1 <= Ru[0];
				MULT1_IN_2 <= 16'd21;

				Ru[0] <= Ru[5];
				Ru[5] <= Ru[4];
				Ru[4] <= Ru[3];
				Ru[3] <= Ru[2];
				Ru[2] <= Ru[1];
				Ru[1] <= Ru[0];
				upsample <= SL1;
			end
			SL1: begin
				Ru[0] <= SRAM_read_data[7:0];
				SRAM_address <= SRAM_address + 16'd1;
				MULT1_IN_1 <= Ru[1];
				MULT1_IN_2 <= 16'd52;
				MULT1_OUT_1 = MULT1_IN_1*MULT1_IN_2;
				ACC <= ACC + MULT1_OUT_1;//21
				Ru[0] <= Ru[5];
				Ru[5] <= Ru[4];
				Ru[4] <= Ru[3];
				Ru[3] <= Ru[2];
				Ru[2] <= Ru[1];
				Ru[1] <= Ru[0];
				upsample <= SL2;

			end
			
			SL2: begin
				Ru[0] <= SRAM_read_data[15:8];
				MULT1_IN_1 <= Ru[2];
				MULT1_IN_2 <= 16'd159;
				MULT1_OUT_1 = MULT1_IN_1*MULT1_IN_2;
				ACC <= ACC - MULT1_OUT_1;//52
				Ru[0] <= Ru[5];
				Ru[5] <= Ru[4];
				Ru[4] <= Ru[3];
				Ru[3] <= Ru[2];
				Ru[2] <= Ru[1];
				Ru[1] <= Ru[0];
				upsample <= SL3;		
			end

			SL3: begin
				Ru[0] <= SRAM_read_data[7:0];
				SRAM_address <= SRAM_address + 16'd1;
				MULT1_IN_1 <= Ru[2];
				MULT1_IN_2 <= 16'd159;
				MULT1_OUT_1 = MULT1_IN_1*MULT1_IN_2;
				ACC <= ACC + MULT1_OUT_1;//159
				Ru[0] <= Ru[5];
				Ru[5] <= Ru[4];
				Ru[4] <= Ru[3];
				Ru[3] <= Ru[2];
				Ru[2] <= Ru[1];
				Ru[1] <= Ru[0];
				upsample <= SL4;
			end
			
			SL4: begin
				Ru[0] <= SRAM_read_data[15:8];
				MULT1_IN_1 <= Ru[3];
				MULT1_IN_2 <= 16'd52;
				MULT1_OUT_1 = MULT1_IN_1*MULT1_IN_2;
				ACC <= ACC + MULT1_OUT_1;//159
				Ru[0] <= Ru[5];
				Ru[5] <= Ru[4];
				Ru[4] <= Ru[3];
				Ru[3] <= Ru[2];
				Ru[2] <= Ru[1];
				Ru[1] <= Ru[0];
				upsample <= SL5;		
			end
		
			SL5: begin
				Ru[0] <= SRAM_read_data[7:0];
				SRAM_address <= 16'd57600;
				MULT1_IN_1 <= Ru[4];
				MULT1_IN_2 <= 16'd21;
				MULT1_OUT_1 = MULT1_IN_1*MULT1_IN_2;
				ACC <= ACC - MULT1_OUT_1;//52
				Ru[0] <= Ru[5];
				Ru[5] <= Ru[4];
				Ru[4] <= Ru[3];
				Ru[3] <= Ru[2];
				Ru[2] <= Ru[1];
				Ru[1] <= Ru[0];
				upsample <= SL6;

				end
			SLV: begin
				Ru[0] = SRAM_read_data[15:8];
				MULT1_IN_1 <= Rv[0];
				MULT1_IN_2 <= 16'd21;
				MULT1_OUT_1 = MULT1_IN_1*MULT1_IN_2;
				ACC <= ACC - MULT1_OUT_1;//21
				Ru[0] <= Ru[5];
				Ru[5] <= Ru[4];
				Ru[4] <= Ru[3];
				Ru[3] <= Ru[2];
				Ru[2] <= Ru[1];
				Ru[1] <= Ru[0];
				upsample <= SL1;

				end
			
			SL6: begin
				Rv[0] <= SRAM_read_data[7:0];
				MULT1_IN_1 <= Rv[1];
				MULT1_IN_2 <= 16'd52;
				MULT1_OUT_1 = MULT1_IN_1*MULT1_IN_2;
				ACC <= ACC + MULT1_OUT_1;//21
				Rv[0] <= Ru[5];
				Rv[5] <= Ru[4];
				Rv[4] <= Rv[3];
				Rv[3] <= Rv[2];
				Rv[2] <= Rv[1];
				Rv[1] <= Rv[0];
				upsample <= SL7;		

				end
			
			SL7: begin
				Rv[0] <= SRAM_read_data[7:0];
				SRAM_address <= SRAM_address + 16'd1;
				MULT1_IN_1 <= Rv[2];
				MULT1_IN_2 <= 16'd159;
				MULT1_OUT_1 = MULT1_IN_1*MULT1_IN_2;
				ACC <= ACC - MULT1_OUT_1;//52
				Rv[0] <= Ru[5];
				Rv[5] <= Ru[4];
				Rv[4] <= Rv[3];
				Rv[3] <= Rv[2];
				Rv[2] <= Rv[1];
				Rv[1] <= Rv[0];
				upsample <= SL8;
		
			end
			
			SL8: begin
				Rv[0] <= SRAM_read_data[15:8];
				MULT1_IN_1 <= Rv[2];
				MULT1_IN_2 <= 16'd159;
				MULT1_OUT_1 = MULT1_IN_1*MULT1_IN_2;
				ACC <= ACC + MULT1_OUT_1;//159
				Rv[0] <= Ru[5];
				Rv[5] <= Ru[4];
				Rv[4] <= Rv[3];
				Rv[3] <= Rv[2];
				Rv[2] <= Rv[1];
				Rv[1] <= Rv[0];		
				upsample <= SL9;		

			end

			SL9: begin
				Rv[0] <= SRAM_read_data[7:0];
				SRAM_address <= SRAM_address + 16'd1;
				MULT1_IN_1 <= Rv[3];
				MULT1_IN_2 <= 16'd52;
				MULT1_OUT_1 = MULT1_IN_1*MULT1_IN_2;
				ACC <= ACC + MULT1_OUT_1;//159
				Rv[0] <= Ru[5];
				Rv[5] <= Ru[4];
				Rv[4] <= Rv[3];
				Rv[3] <= Rv[2];
				Rv[2] <= Rv[1];
				Rv[1] <= Rv[0];			
				upsample <= SL10;
			end
			
			SL10: begin
				Rv[0] <= SRAM_read_data[15:8];
				MULT1_IN_1 <= Rv[4];
				MULT1_IN_2 <= 16'd21;
				MULT1_OUT_1 = MULT1_IN_1*MULT1_IN_2;
				ACC <= ACC + MULT1_OUT_1;//52
				Rv[0] <= Ru[5];
				Rv[5] <= Ru[4];
				Rv[4] <= Rv[3];
				Rv[3] <= Rv[2];
				Rv[2] <= Rv[1];
				Rv[1] <= Rv[0];	
		
				upsample <= SL11;		
			end
		
			SL11: begin
				Rv[0] <= SRAM_read_data[7:0];
				MULT1_OUT_1 = MULT1_IN_1*MULT1_IN_2;
				ACC <= ACC + MULT1_OUT_1;//52
				Rv[0] <= Ru[5];
				Rv[5] <= Ru[4];
				Rv[4] <= Rv[3];
				Rv[3] <= Rv[2];
				Rv[2] <= Rv[1];
				Rv[1] <= Rv[0];			
				upsample <= SL12;
			end
			
			
			
					
		default: upsample <= SL0;

		endcase
	end
end

// for this design we assume that the RGB data starts at location 0 in the external SRAM
// if the memory layout is different, this value should be adjusted 
// to match the starting address of the raw RGB data segment


// 7 segment displays
convert_hex_to_seven_segment unit7 (
	.hex_value(SRAM_read_data[15:12]), 
	.converted_value(value_7_segment[7])
);

convert_hex_to_seven_segment unit6 (
	.hex_value(SRAM_read_data[11:8]), 
	.converted_value(value_7_segment[6])
);

convert_hex_to_seven_segment unit5 (
	.hex_value(SRAM_read_data[7:4]), 
	.converted_value(value_7_segment[5])
);

convert_hex_to_seven_segment unit4 (
	.hex_value(SRAM_read_data[3:0]), 
	.converted_value(value_7_segment[4])
);

convert_hex_to_seven_segment unit3 (
	.hex_value({2'b00, SRAM_address[17:16]}), 
	.converted_value(value_7_segment[3])
);

convert_hex_to_seven_segment unit2 (
	.hex_value(SRAM_address[15:12]), 
	.converted_value(value_7_segment[2])
);

convert_hex_to_seven_segment unit1 (
	.hex_value(SRAM_address[11:8]), 
	.converted_value(value_7_segment[1])
);

convert_hex_to_seven_segment unit0 (
	.hex_value(SRAM_address[7:4]), 
	.converted_value(value_7_segment[0])
);

assign   
   SEVEN_SEGMENT_N_O[0] = value_7_segment[0],
   SEVEN_SEGMENT_N_O[1] = value_7_segment[1],
   SEVEN_SEGMENT_N_O[2] = value_7_segment[2],
   SEVEN_SEGMENT_N_O[3] = value_7_segment[3],
   SEVEN_SEGMENT_N_O[4] = value_7_segment[4],
   SEVEN_SEGMENT_N_O[5] = value_7_segment[5],
   SEVEN_SEGMENT_N_O[6] = value_7_segment[6],
   SEVEN_SEGMENT_N_O[7] = value_7_segment[7];

assign LED_GREEN_O = {resetn, VGA_enable, ~SRAM_we_n, Frame_error, UART_rx_initialize, PB_pushed};

endmodule
